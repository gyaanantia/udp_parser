`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam PCAP_IN_NAME = "../test.pcap";
localparam TXT_OUT_NAME = "../output.txt";
localparam TXT_CMP_NAME = "../test_output.txt";
localparam PCAP_FILE_HEADER_SIZE = 24;
localparam PCAP_PACKET_HEADER_SIZE = 16;

localparam CLOCK_PERIOD = 10;

`endif
